// Main Module
module led_driver(
    input logic reset,
    input logic scl,
    inout wire  sda,
    output logic [3:0] leds
);

// Power-on-Reset

// oscillator

// led_controller

// i2c instantiation

endmodule