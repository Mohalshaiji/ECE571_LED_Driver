// Main Module
module led_driver(
    input logic reset,
    input logic scl,
    inout wire  sda,
    output logic [3:0] leds
);

// TODO: make reset active the same globally!

// TODO: power on reset? or some sort of self reset

endmodule